library verilog;
use verilog.vl_types.all;
entity testMreg is
end testMreg;
