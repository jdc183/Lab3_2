library verilog;
use verilog.vl_types.all;
entity testAreg is
end testAreg;
